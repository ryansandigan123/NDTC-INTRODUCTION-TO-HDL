LIBRARY ieee;
Use ieee.std_logic_1164.all;

ENTITY LAB2_PART1 IS

port(
S1 :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
S2 : IN STD_LOGIC_VECTOR(7 DOWNTO 4);
HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) 
);
END LAB2_PART1;

ARCHITECTURE Behavior OF LAB2_PART1 IS
BEGIN

HEX0 <= "1000000" WHEN S1 = "0000"else
        "1111001" WHEN S1 = "0001"else
		  "0100100" WHEN S1 = "0010"else
		  "0110000" WHEN S1 = "0011"else
		  "0011001" WHEN S1 = "0100"else
		  "0010010" WHEN S1 = "0101"else
		  "0000010" WHEN S1 = "0110"else
		  "1011000" WHEN S1 = "0111"else
		  "0000000" WHEN S1 = "1000"else
		  "0011000" WHEN S1 = "1001"else
		  "1111111";
		  
HEX1 <= "1000000" WHEN S2 = "0000"else
        "1111001" WHEN S2 = "0001"else
		  "0100100" WHEN S2 = "0010"else
		  "0110000" WHEN S2 = "0011"else
		  "0011001" WHEN S2 = "0100"else
		  "0010010" WHEN S2 = "0101"else
		  "0000010" WHEN S2 = "0110"else
		  "1011000" WHEN S2 = "0111"else
		  "0000000" WHEN S2 = "1000"else
		  "0011000" WHEN S2 = "1001"else
		  "1111111";
		  
HEX2 <= "1111111";
HEX3 <= "1111111";	  

END behavior;
